library verilog;
use verilog.vl_types.all;
entity decoder_2x4_vlg_check_tst is
    port(
        O0              : in     vl_logic;
        O1              : in     vl_logic;
        O2              : in     vl_logic;
        O3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decoder_2x4_vlg_check_tst;
